module SimpleWire( input in, output out );
	
	assign out = in;
	
endmodule